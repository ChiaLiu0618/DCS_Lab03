`define CYCLE_TIME 10.0 // Cycle time in nanoseconds
`define PAT_NUM 1000    // Number of patterns
`define MAX_LATENCY 100 // Max latency for each pattern
`define OUT_NUM 1       // The number of output for each pattern
`define SEED 5487       // Random Seed

module PATTERN (
    clk,
    rst_n,
    credit_valid,
    credit,
    price_valid,
    price,
    out_valid,
    out_data
);


`protected
[b64LGZN6a))XR?4N#]>[L&5T=WM^>FMAI<Nc>IPU4<fZ7dM=LWS/),YGIdM__HO
d73<b[a[+X>+L;cGbL<NC:#Z.M8Y]P5];Gc[R8R,(UDGggBH96\b3F_[GW-4_RdA
/+dYIdI5f_#U+\aM8XL3EIGa0ZcA)@FMbaE]@>7CAO8F0,M16E>O:Yd-SPP7U8[V
5DV/QZOSd&(.U(W]75Y+X17Rbe4(d/,FKd(>5KDMg_VZC>^ce@Oe6F3]P74/)YS;
MME_R><_Q.Ic8,UD.8DX--<V]876674,T2(V@7&_6OZ8>;[82B7_42:a9]Cc@516
TGR>C)V=-CNc0$
`endprotected
output reg       clk;
output reg       rst_n;
output reg       credit_valid;
output reg [7:0] credit;
output reg       price_valid;
output reg [5:0] price;


`protected
aV=:]@9P5UP1a[)RcC5\B#N8?/cQ6J8T0;XPZ#P08GR)<+QZ)AdO/)=Z)DYgJ8QL
J@:>\O;b\4WaE2_#O)-A76,C94^6&2.c:$
`endprotected
input        out_valid;
input [8:0]  out_data;


`protected
)717)_<@2PZGCEB.FMaZ:IW.IOAP4A3d73NT,2^=)V(&WE5D?DbW3)X9II=2e:\a
/6=PP.+e5Y-.+]Dg\UQGeP&]7F5^CJ1O<]8W9N(VP^R8=<JQ347M?O0WE8#b-#.<
Yf-(PF<:[&BC:gL:(]INRUP.&^Y5JUVS)3/d)aM>1)&L=1G21N-f#]L)SfQ,>P.X
c2NIf0T;.@WXJ=,WA]^.,C&/f=QdXaJ,c98HPRJ@YL,+))D<-CILOAO6LW>3b=Y#
)1.)F-)TC9,B?8X-X\;HgM,F^OY;Ig<6OBQ>XM?)YBe^VG:\E+?eeN;;OS4KGN=2
0U()[c;:WY@[Fa:Q\gCT8</C3G8+5G:NB#2S#NK<f=2IS3^c?2FGaOD</H&-PJ+a
#ONYd_@KY;74;fNe:eB#[AdO6]))X,X948HGaT7ITH>Z6LX-QD#QRL3Q(PfVX8J]
Q5H\]gJ9dK+R35W_SB2]f#-JMV>N)da-TP=L4-V^H(eQ0S10Y(AK.CfFK_[D:-0a
?cZ(;+^2b6@[V?bG5EVB,Kg]K?HR>_PE2AG@]K_TH&f<b3A62,+OZ[7gA]8#./V?
SG&RLAQ\gM=?AceWYK_.Q4(2<#G<eF/#^TdU;g8&?5=#.\>O=JS<SZ3J?Mc6:91I
c>XP@&M(Q<LCXN+O:dQ5:7IB:-[Y>/W]g2&_^X&(0dZVR:9XW448[\INS/WD?FLa
+c4A16@b:aDSQ8+F\d0GRH:(D(g<1<9DWVR2AL-A#3UD):(#W>L3<W+>d])6Z0C,
])ZPB]VReZJ/<WOQ4&&3^aFP]G3R[1?<IfR<e)&H_R6[f8TdVZ3bN]d>6N,V^8PZ
_</g2Y&@8Be.1[K^E[2e#Q[CORX3,_=KN)SJgGRH3;[:PR7cOgII]S2b25fE<d.3
2N2,R<.9]<5L(M[^#^Tg<TL,Gf:gABJ@g/bFc/46/[A+]5M4(e[>6OcgQc>1\U>9
7bSS\3E;?9BW/eNd)HDAF\L/1b&[)9C8VFb4E4(3\YV;&5B44++;Q\g@#HHO^)6?
d;6XSVQL9CfGRX-_(:XDdRXXNK.J1@/3e.Q4VP:0a:^L-()D][SQPFL3AB.WE6>1
?MF]B,8c.>M)1d+E)7+<L3a)V;O?@[GAY=cCSILGM-0X>9QGVHD;(2gXO:DbdIVL
[H[+S^GY;W+f5;Ic.N/<.Y^E0WZ\+b43KIC@\)>/1(#.823=KKSC-58/0D):eKG[
)64GMYUU)[XLFE;5ON<V?>#fG=JN@U]f9A_[78g?/5F7aS+:SQFCCf:M#^T_f@Z1
Q]GYe+7,&S@D1B9a^-(JX0R7dR)d=_7=)#Q[PT1L7:C=cdA@\#(eM-7(bQ&0RKEV
TBF0HdN\?[d2K>DUMdS?#_2gC/0(SMKBPL_HFT:[g8UJ28)P\W+I76bbVIFNZ2,0
]YQ28JHf:OC).4g)=74.?QKa<O14Xdc>3T^a5?da>DWDVP=YG&/7D=QUDf/g2//^
[MaRNL8@9dI)#RBdVY6)e=G_2W+XaZSB:D2CCTMOcP?:>fb9T_2K7WI12L,?UB;2
f0Y7fffSZ2?A9Pf(5+Yc/&Y5Q^V:K6GK1HNZd5P?:@>ga6D4P4HfROe.,IY\S\>;
DVEa+@&Xb0JgXgZa\V?-#2.T\g4H6?;-d?YO@.OV<[:HY4KRaX=[c_S1HX>C87Le
a3.?7DNZ&5;\5/L\_\(Zc6AE+gFI/=-T4MLK)P@8C,\F+:0(#NBTVecH07(8?#Bf
<gR-IfJ&.S-g(&L=PU_E8U,aYg(;#U[@GLYeJgBdQ34F;Z]OQFa2<[b,>;ZLT5U1
INPb7;bcB,R^=[\1)Q\(8:?ENf]Q1&X.Ia_NE:ed3.=@F>K>bWgKRa>QaY2V#\]d
QS_D]#N8cPA#QQMf^8JZ5NEC3J9JZN2P8fH1FAdE,U\cMD5BI9\ILTK)OSZ)OJ[C
H_ZN:Fb<CA=R6c.XT<.N]JXPL/RZZcC8?-4^#_d/e2SACVEMLA,b-<V&E:NS1210
)5Q\F=LX1AYY1(_g.O?;E4\#SZ4A;(:D=D,.,JN,RVVb_?L<(8IQb][=B^KM\#g-
L#A[X;fI?#7H<,@ZLOC[1[#9F3=E4EI)=S4bJY(X)IZ8J0W+>]/JK0N-QZ8D6DI>
+LVN#dX1]NffUN:X4U12KDQW<4,F.b>4-0?X/e5R2U[&R6/RD+##>#CY;a)H_RZ\
6d=f\T;57?:HKVdKE036_JE9_80U+6FGeGfELSZFR>Na^c9?AJJJeH<UU7#-1T1c
5&SDg+8dT8(;6d-[fPN,<GJKYg/gc:4^Pe2TDWdG3@BB1.f8PBa:dW5MF@GM9KBB
e.PYB_@SRcBc[gdN4eMY_0XeS>[==J^@^XFf2a5V)\DXZd3C>=A=@2O_5Vb54,([
_&8:<R>c7F4=F8c83dP-E;VG87D=f67b]0],R6UYNIHNfd4,C@>42:[d+agU^&Q(
X/>OK\EHM_J7F0DM]MdcDW2CFHORH.KM7LI7#FX.HI\_5UTRK/.^?ECPTEa_55ND
Tb96-7eR>MF_FDVT\?)^>B;61O7&/(Z5V2f6_-I#aA=gXf#0<[ILG457O^L-8X+M
@HIff7Ag>8H=99/F/G&AL5S.+/g4-U9YSWg\4CXSe_I7F]fLd/9@KAc5&6VNUW8?
OY=4SAKK\IWVfCM6_ade\<P3Y&d4<45QEEO8gNC&aF\H0bI&IP@bRXg-Ld3c/AXY
A\fJWR[F__].:BcRcL[\0\QR&;f=&S(K=@D<X:8WB4H1_:;b]L]Q^>/JdY](<4b2
OP@&>:6<4NP\HQLUKG7->TZ&LLI]Jc;=dJ\FMfO.BfYP;U2WRFGE7c8>U3g9HRC=
b9>FfPNa.g+)8P<W:CM289HHU&\5WV1Y\S(b#O@a;LbX(UdK]9SFPa2XHc\DadV1
=c9^7A>5DBHA8#9AV0KO^#8UOJcDDIfJf\,YFKHK@J-])K@_.0IUg.U#JcQR@T)X
.Y@\MUGA-dN)g?SWD1?,C]?2\6NPG6=/U8K]#SH-MfAP^Og7H,5aS1GPcGg9V/1H
_H6A=[UXL4BLN8UD?cV4PNNBA4;Y=+[P_+]Z4FCcDE>&;-J5BQY8eb;X90BK.2/g
;<BWLgI4CfVTP28&5YMI@B]_;\0g\^d5(F#9QIFgcC_Z@)S-F5914b6Z4MD45#-g
MQ(QdIML)73(:.N:NE_S;]H/7_@bL]^,937NUNYc)24a]UZ2/U\(1)+X=91\1He/
,Bd=L3+]b8BC2SG/:SXbaBKcHEP3NW=.BS[@AUe)L_f(EgfDCc9#+8V7/I2=XD75
2.1MGTc3\dS.bV^=5L0YTC=?EMEQ99#b5\CGg(TYT9c,3d8I3fg)_NUN)#;[[)#a
T<,=ZD(.9RH)VgS?>LF@5<<;HD7a#.\C)Fg3AKbZ@93[XIB(3O\B?;/BUg#0:5_V
94Q@UWacE&_7JT]5>[/=0HPSZ5@ga]]MN1CBGIO,XVb)M@^3Re4Vf:)G^;JOU.]5
9).N/^BV(&_HJc-3I((/IZ;N^R,6>GO?[,(2b1BTY)T,N9246fd)0^e1&#C3#@d4
I>gU2PfRfaefHLIO3/V<bGRKW7W2;eF-+NHL\(1d&.\XNeLV+>CB]MQS_87\SAeF
H[7K.CZZ1Q,+I@YIC7XRKGW.\d&E7ZSa8dMK-K\F:>33AdWX#=>N^1HU)#PU9_U#
FLaB]M:=EF)[E;3.&5d5V4BgJ6+eR[bGO4JfF5d;?EY./e4f6.\G7GPE@(82ISB<
()eB8_(>#cO&Y_aaTV^DREeSHE0][^^agP/c9AYWdEAb\^WR3E2/C.?\BR/e+/YP
PNYVSC0O:,>[YJY_]U:23;ggK(OUca?OGD25\[1c\P_7-&aN4?7g9-,NKT36\6BD
fDU\(HV2g8&@:E:5F@^@USe66@0QTAW;:N&R)&O-fBR947HA^dPH66=CU-2>R^U7
H0G=[?:#EVR#8\4.^.T+>8e=8XHDVOKC##8GQEMcZI5,#XPd:3gF^McP0Z,g9JBd
Tdd646>TaB8&aN?E4T(=1g\,PE?(g-6;&=W=gd>TO,Sc3fWOaH9XI#NIGI0#L9fS
6<O0<=VNM^AXXM9Zb.8d46;a_\C:#FcadX#3^Q^K/-YAW7U_43HBbeGJ@?]K\I2@
TFZ5F;S7R1b.F7,RC,U]EaPfY:.5F:LfG7R62K+21,>8dE(([53/IXQ^,4Z?2,]U
<e#B<>)cAZJX+_[7__-05#:\2K._2@P6=B<8M?a0B+K<g<DK5X.]U?7L/ENAgcYZ
d35FS0^RKd&.c<);D+TPV9#:b^Vb1/)5R.JT0bT+^B[^@A_@^\_<7RL^.V;W][&4
54.0dgVH;^-T_UM;Xe.3.S9_K[7b3B,HMUY[9[LK[77(6@cWYK^[WOO<Gd367AE)
,/A_&KME2=Lb(.d)<2:W/d3G:RfYO0d?HF5_\@PN;a=UF5FPUVDANaaT&P(Rgd^@
d,B/L@dDf1g)\TJUK/1a@K,bP2Q3TJ&=\FQGJ>e/3Na\/&.e:&Fd=AgN+HPM^5AE
[V68cILUA29M]6O<X:#TPJ6DV03cO6f82394g=0(d0Ge(13@SL=eL6,4b+1S9@US
](U2E9SXdGfW1C5gNbOK1M<7_^B+TEN.;E&AHaDWa/MUYYb7AC80=@\.cOXf.(T(
?E;>E>>G<U)(P,bG?NeE[2;Z?=KL>R]Z1GK_L5ca)SSM95O6_U=<PF5FWEd:OGWW
M^6g=G6K#baL7W5:DQH4dZ8>a;,^90=T6-#SY=_SFOMVEDQ3+ZT29cEcLg+d0[;/
DQ8;>5g8(\ISRBU]A,[RL/dV[PVNYg-2Y/(4KfG+)O/g-f=-180S)(8S_GR?&Ecb
D:fVY8dRS9(SZ:gXXA@ZQ6a-U;3=JI6c3@+f&J8<8_T2-SQK&b_EZY(46J;?84Jb
F5DJ)N#gTSaZCTc&dB+@5GZFa5QJBN&Q0DS_>#T787@NX(XEIM#gB(2_a(E&C2Q.
Rcd@J+S>?ZSdQ_;cKHK5Z3D7G#TKg4>I.-ZP3@_&IK@F>+g9_QQ+WO9\Kb77G::Q
E=)8N3Y]X&4KEK2H/bS?W\GZ+d9O1(I/VS]HSbPS5QI-9I<XCFF#OdKe:^e,^@AF
fTUgBS<3FYXQ4I-I>E[=#GYeYK/#1LWW>Q.[?\g\7B[X@4PAN2e,4946TC=K#_(#
Y9.?<RV9NG:5Y3bDCaB-O>Q35:edB8O^A^Y<OQ<\4f1/N[#L3B6f/PTeJDO?-FgU
@6^69/D8g[88[fe(<a[0[S(A+R>VGC4?Mg__#WGXYc\d_c4ULNDNK??1745W+0Z+
Z<G6f;f\PHacOgge@2HF+WO-0@8EJKZQ<D5=N-/@E[fU+;L1gG=83QaWWD^55P.#
/eQE7eDU-T^L)6:8D&df_(fFBJ3M\aKKUIMOOWTM):3GHY9+D17+fLB:#FCaX[SY
^Y_3,/fJbdVZJG<6L9b6&\<J>1L.<AReeFIMPaW.G-5L2CG@2H4E3dA9DRZ3g02<
PaEASg+KWe:EC.51?W6HH8T@IK<UX0>&A,6Z46J81ab\JC6g9O(_:b=;)6-O&F>8
WR.R6K(Bb)V]II7bR:T)0KW(a-2_G)RU6AeQF^5E]@+^OY8+UXg^VV#)-6b]541,
AS?G@M4WV+DD_+W).O[X[;8L#;O&ARQSa&T>-^egB;IbR)(#)0=C,1f[QEEa6J_W
=7(7Me_TYKdWN:NCE)6AIOgL?2K?(YP=0Uc&e<72c#9<bZ5IZQVVPccHT[+IX76Y
MDH+=3[db>&CT(R<0VBNDCg@:A,K8--/P3+eJNQ]Y;MP-/+Q@>):)STS2QJ\VA)>
GV)ZDZZ/E2&IM]^>c8+0[.33+P2NgFQC.G&TcDU4b[\=KGJ99H7=;KPNOEGJSQ=:
>6\b4gS.5IT@3TL0T<<RW5-D03.;BcOW6>4[0,YYB,#^G4+IESKV6Y\aDRQBAGXJ
[<8ff[[f,^WLL2+U7@bG\/X>8;IP?RabfP6+80J?d;M/RfQ0+)Q@HXV<a8G6#E>.
g:LJ9Y=,_;;L&^bE?P3X(HAM4F/C4CWLN7e^0MVBB@8#EG@9BY/;C/OP1KH8E6^,
,99I=^N&YF&^[fV;eD)ggY.DC/46:=(Cb87C@4HEcc3gG?29DV/@+#=DLANW@NU2
0W1,5OO]K9TR6Pa7X8S&HD1g\Ag+.BBH;3Z1/86IZY(+DW-XLRBMc7Ta2W/^0A24
L]_6b+/VXP_UU4F<_=fEM1NWJ&V+@@]\>65\VCC1#(66SA)^>I4,9M&:Kc/d2Z1]
-^W>bH[._]/.556JX]=8N^\/JN/cS]Jg_+XEC:<?_[HB2bB.9>1.K9GP\HRKXAIC
[52L@TV(W:?XQO-TB_QZgCU9<(MV5K6I>F[VdB>S^Cd?HKe#A2Rb9,9VLPb>5J,a
Wbf>NF9;V4WaRee^Lg[GL]9RZROD_4dTU\:#:<c1bPRGB8V2e2cNF=YEUEQcQafb
D-GcY[J+HAGa7g4&?e#+<<Sb)5K.@&<>=XW>^VU6HJB).Q^7#L^@J3#9;_,^CXIJ
O7&P644>c-IQ6)AH\04b46,X_;MHNN;&KIFEOc0?EC@I1R#D46MX7/:C[TEEO0eV
=V?T\O@]We.&+#@P3T(:8GU6]OFAL&A7bPV_I8.d/_c:@=JQ2F:I?>D4NE;,F75>
H67#HedbMAd#T_)DPUJ8ge]1LLW2)Y15:cZbB8X&cc[fbHgSa\WMPY,fNT5M8GID
&AVAANU#eb0SGR3)2VH05NNBC-A23f[X[X+#f^E=,5((@45]LY4#.TJ//g9KDNRE
7:WSS3?8b7Q6;(4\CV._Z;X?FL=GK;X-WLJ73X1UUTAZ<_Hf08P&9KB@_4g3&6g;
GAZ)DF)]2.>G:6Ge6^b:0B#;2P:X\<\]NKQ;,)X^F?V:Q5&W<_0:2UF1NEeMa37b
U6T@EFd0QLF[?M]?H&+FX0<+O[H/W8bE#=WWI9JK.D:SYJ,PD[D(RKCW@7b3H0V=
3?bL2IXC_UB=+b9A7/]6bZa3P@1-Va#[PG42R](Y_R1_,P;?d@>@(A[<X6.5feR,
dC#6E\4>J;Nb[RcWK.Z_Y:Y26TK89V<4):6IIO9I)22XYLd8Z?4Y&>5^S]aWg3c5
+_R_NA;1,+N:J3FT:CM[CEJ9>7,8eNd3<>6UGP:F:P_U#ZZgIcg.^F3^,L,=fe4_
eGF]9K03Ae@?IKW<Q6\KOKfUZ=R6-ZT.LZD8#^R7S50Ma(@?fHB=^VTNL<^+Y;N)
DK]aKDgFE#?=Ta2[301Y3fH[ce,>B+Z;J8F1VPSRNPKQOO-VQ3.ZD.QgeIPDP8Hf
#8@JIbCU4L=LG55N^#R)8<E[.DBGFT>FXf(D)bS&N,a7&5SMaP3EZdH-,)\eM7\B
^?:9HO##W/HHG75e1,K+>>a[-?SM<[TRB=#U8_:N7ddJE2Y,8PGD#>RBLTOA#80&
_<aB5#9N1e0@\aI&>3///<^(;bW>A2e9;-AQ:e8V(5db]3f9YdG)b2T3V1D(_>-Z
db@+?ZISM+_c5eJ@YK.DFCb7MGAZLD#[,\1=Vg5JfGHJ.+0gcf@FN;+O^[LO8-AG
a,_A^E8.UH94GY;1UQU]9(/.)R2A>Y:>0<V;@=Q_&O/=9Of8O?:G0>Ue>^F_L>B9
S?K\JOPM-Tb7QJWY[A[=SDf?H(bONgP.d[@W:Vb5.aV)#M33LBX:DS,MP>5S8LaB
:e>U:;@TJ8)#TCSDe&3RV,F#Q1:>fIW#TagALD]D6F>>1aWgLRgVXX^]T#\]]ZfG
QIC0[EfQJ8G==.H[XG^EXONTYH[V_Ve&&Y0GY#)IF[.YUO<-JD.b](D-JOJF?-M2
RPB.c3PHZA4\;]fNH,AH&HKQU#AP/5BS6?F2EBP_JLZ;@#>F/b-B+DJ.EfP[aC3g
a)XW&_S1I.eSD/-/0?U/_?.^=#D\ebe-I3d(HW9W)CEAR+H64QA7Wc0<3-\M-3RY
OL]I<Y01CdTM3B7Y):\<gV28D:UN?3R;gN&e5MKR#Md?;V6NL_0&Ob7B@B8[VV7f
_=QP.B,cSb_5M.LQb&BeP,,fE9f_3cLC358I,^9_PWI/D>A@(OE1JdU#QPM#0T2S
ZPNZ;=aM<W9eCL0[:FF]7d.A#&c(1.I=:]T9?,,[+1SfLe@^b6d#KN#a=H;)\[RE
=G]+ecS:b]3e,IHfbe7WG_[If-)fdB]g@c08/NPT0d/W(+EGaBN]O6+T/eRB<f:8
J.DE<X1MX5ZZ9,Z<cK..e-M0.EPXXE^IFg1]1Lb5^&I5]6==7@1JdbRK;L),_EW8
\b-NJEHg<;L>^R)_M@GV4,FW?W<+_3C+D7VD1@4BW#RAg6@S0:.T5\@\X0&6V<dZ
V@V.D\7LGYd6<&(3M\M\Z=EC3.;>E46.F@&9I5Ie(fcgD+.(8Q+[<<RQ<K<V<Y=)
_UQ0S=b?9K7\Pe+@>FCC)&gMUcO>UO7>>,L3Y.+=KG)BC=JAXJ+,874,Ye<>1b;L
P:/eBXg06Q,ZNc38Q]QJfEdM3S.G2WRHS>MFHE:6&(D_Pd1HRg>WEDIffX.^I95e
_]NR1QO]2]WD)T?BOIE:aOBQMB;A>]-)BeR(+>O@3I<QV\eY;\MW(@H@-F7C.Q6)
JAI[&KeT8IS+DZ,Xf<2+IOe)QXdH@CO)<b9J.1\2ZP5C98.YD-&/HQG92,g#2I:g
FP6[f8+^_,\+=d3XE#CRFe<3MeTRK()F5g),OX,b?]B:)<bXQJUSdEQ<T;U7VHTO
?PbT=Z9^g]I,a/JAfYK459Q#Z]A?K^&OOFGZ=e>21IeHUMg)YX#:g/>gL6=C5.4A
C5R>2[M?UJgNC#)9cB6U#K.]U<?E?W)[ED.]6fTc@fA(g<<cPFL(e^BbdeM?,&f,
)?a.K6]VK19D12_aYf1<_\9Q?]NPd7:-_<6SU2Z6RM0C]^2X^Id;_b#/]QI4PVPH
I4USN)&;JZ?^TX\3aX^:@/Tc1+]UPee->(IPfXYQBa(5GgTaQZ1Z^>9cef[^)]d,
4N?XFa4?46J0>GWK_-B&^-;H,c3-0L\?C-g\:<1X^4-W[8-Lc@49DaAQQ2+PAU][
adS(NJ_F.[&+d;-=PJb,\@Mf5FW18:/0ObKQK23]cV#L6HEQGTF;3/=P9\-KA^5g
?gN=XY=Q<@96:I,.,HcXa:g[./?b[1gV[c7MW85&R(Bb4g>:Nfd,BI3@a<.ba7Fa
d(7TS,:_WS+31+b;HMA\;N_M-]&a\S08.,B>0W,(Db=)c56C)gaC>(9H_7gJ]BIc
Z@)Me:W7RI#TPC_Rb.9BX5d5?X;S:HaMY<-bOeVOQ61T)a.W?JOH)(?dbF#S)c3#
JNXA@]I,TF_Y^9c9beZ#L&Ad,.8S\65=MY==9E(2D1VeJ:DB]\ITa3<W[[T59#TP
X(F2Y(@=aNFNCK+T6PJ4EICT?(XX2.V_S8dfeKP.>MMHQe&I3@+a/?R]J?72QSf8
EE+Bf\>+dNaVXHLf,;e7NR^5<S(aBJJ)?PQfdA=L#,ORJ9E)BRNg0(]+WE91EPB<
B86FD.-BV\FMEA,Q-cAb<QR>eHT&+X\QdO>(>,EUSAJ&=(YYH:\U)@E=&aBZ-./&
]F@f//M56Z3>-Nb[FL[Z4Pab22.F?O&cDT.U=/afMD/eaSd9cU8-NF=G[01[=-Vg
C]I0VbKb&9B/X+<E=XPa1O@)5(/Z\Y68:7VB@R/7QJ8.AJ1bbG9)d4+cK@>YUY-G
YYAebAT>\Z\g0__T1MM5C5ReUgD5bD1:;KL_/:4f7f,+a]]GJ_C7gXc-KSMHe;g<
E;N99^0J28;bD;/dNP=R-?_PbfE&D&[-0H2(+,Kb1?(^;<a;3_G^X8VYZFFf623T
SXA3]a+[SdPaEaDVZcd4aKcB<-Y8bTNcJDI?P0UUI#X?f^>WPK3UH5@R5W2cAXDP
Zb>>=LA3-[681ceLQU6Je\G;N?,Zb0UWJN\JK+IEYYT28_;Q1RUM#>3d=/<QE<O>
UU9,HCg[_TUD=)d5P[?E9-&aXg[3JW?L.BdNHX2gK@],POTO?_g#:bE/eR9f6[I)
ZPWUW([,Y^8Y#.73W]R^.@DJ;N(dZ3TW#R9-PYUDV,=UQDLaZVKH2RA<&=KSU]XH
F\XT/D73D)Vd0LbB9U_N0Y2cE:RKH:T[-:R=fa(V,>PUB_gSO.CSgC6b5IQa;PG0
/O83@M-_Y1C<)^Q&7-f.@9:#<:4b\;KCUPM_LKc#JIe2_J6/K^1@5/RW+F4ZBA<]
0_gD+1O9@&0@T>[-NSNcL8:J.Ye0HLT>GY<L[2W.UE]-WJN,F<=B1+c+J@AT)_M5
R8#dJI@_B]IROXG_)EX_KZ=O&Qg^?Xg:1a@PSE0-A)DVHbZTAY5PAdc+P$
`endprotected
endmodule
